-- <header>
-- Author(s): Kariniux
-- Name: internal/testpy/._tb.vhd
-- Notes:
--      Kariniux 2024-11-21T09:04:48-06:00 pushing-pulling
-- </header>




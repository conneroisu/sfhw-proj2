-- <header>
-- Author(s): aidanfoss, aidanfoss
-- Name: proj/src/TopLevel/EX_MEM_STAGE.vhd
-- Notes:
--      conneroisu 2024-11-11T15:18:36Z Format-and-Header
--      aidanfoss 2024-11-07T09:50:56-06:00 fix
--      aidanfoss 2024-11-07T09:37:43-06:00 create-exmem-stage
-- </header>




-- <header>
-- Author(s): Conner Ohnesorge
-- Name: src_sc/proj/test/tb_instruction_fetch.vhd
-- Notes:
--      Conner Ohnesorge 2024-11-21T11:05:34-06:00 added-old-single-cycle-processor-and-added-documentation-for-the
-- </header>




-- <header>
-- Author(s): Conner Ohnesorge
-- Name: proj/src/TopLevel/Fetch/program_counter.vhd
-- Notes:
--      conneroisu 2024-11-11T15:18:36Z Format-and-Header
--      Conner Ohnesorge 2024-11-07T09:51:12-06:00 progress-on-stage-2
-- </header>




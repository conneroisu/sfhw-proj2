-- <header>
-- Author(s): Kariniux
-- Name: proj/src/LowLevel/._xorg2.vhd
-- Notes:
--      Kariniux 2024-11-21T09:04:48-06:00 pushing-pulling
-- </header>




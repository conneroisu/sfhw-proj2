-- <header>
-- Author(s): connerohnesorge
-- Name: 
-- Notes:
--      connerohnesorge 2024-12-04T17:49:24-06:00 remove-testing-bash-files
-- </header>




-- <header>
-- Author(s): Conner Ohnesorge
-- Name: proj/test/tb_instruction_fetch.vhd
-- Notes:
--      Conner Ohnesorge  <connerohnesorge@localhost.localdomain> change-name-of-instruction_fetch
-- </header>



-- <header>
-- Author(s): 
-- Name: internal/headers/testdata/basic.vhd
-- Notes:
-- </header>


-- <header>
-- Author(s): aidanfoss, aidanfoss
-- Name: proj/src/TopLevel/MEM_WB_STAGE.vhd
-- Notes:
--      conneroisu 2024-11-11T15:18:36Z Format-and-Header
--      aidanfoss 2024-11-07T09:57:02-06:00 fixing-extra-control-signals
--      aidanfoss 2024-11-07T09:50:56-06:00 fix
-- </header>




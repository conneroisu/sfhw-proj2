-- <header>
-- Author(s): Conner Ohnesorge, Conner Ohnesorge
-- Name: proj/src/TopLevel/Control/control.vhd
-- Notes:
--      conneroisu 2024-11-11T15:18:36Z Format-and-Header
--      Conner Ohnesorge 2024-11-07T08:35:18-06:00 run-manual-update-to-header-program-and-run-it
--      Conner Ohnesorge 2024-11-03T11:10:31-06:00 added-a-new-documented-control-unit-for-the-MIPS-processor
-- </header>





-- <header>
-- Author(s): 
-- Name: internal/headers/testdata/golden_basic.vhd
-- Notes:
-- </header>


-- <header>
-- Author(s): Kariniux
-- Name: internal/boilerplate_src/TopLevel/._MIPS_Processor.vhd
-- Notes:
--      Kariniux 2024-11-21T09:04:48-06:00 pushing-pulling
-- </header>




-- <header>
-- Author(s): Conner Ohnesorge, Conner Ohnesorge, aidanfoss
-- Name: proj/src/LowLevel/dffg_n.vhd
-- Notes:
--      conneroisu 2024-11-11T15:18:36Z Format-and-Header
--      Conner Ohnesorge 2024-11-11T08:50:02-06:00 merge-d-flip-flop-into-the-structural-definition
--      Conner Ohnesorge 2024-11-07T09:51:12-06:00 progress-on-stage-2
--      aidanfoss 2024-11-07T09:37:43-06:00 create-exmem-stage
-- </header>




-- <header>
-- Author(s): Conner Ohnesorge, Conner Ohnesorge
-- Name: internal/boilerplate_src/TopLevel/MIPS_Processor.vhd
-- Notes:
--      conneroisu 2024-11-11T15:18:36Z Format-and-Header
--      Conner Ohnesorge 2024-11-07T08:35:18-06:00 run-manual-update-to-header-program-and-run-it
--      Conner Ohnesorge 2024-10-31T09:22:17-05:00 Added-init-files
-- </header>




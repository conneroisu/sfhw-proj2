
-- <header>
-- Author(s): Conner Ohnesorge <<conneroisu@outlook.com>>
-- Name: proj/src/TopLevel/Control/control.vhd
-- Notes:
-- 	Conner Ohnesorge 2024-11-03T11:10:31-06:00 added-a-new-documented-control-unit-for-the-MIPS-processor
-- </header>

